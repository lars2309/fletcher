-- Copyright 2018 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.

-- This file was automatically generated by FletchGen. Modify this file
-- at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;

library work;
use work.Arrow.all;
use work.Columns.all;
use work.Interconnect.all;
use work.Wrapper.all;

entity fletcher_wrapper is
  generic(
    BUS_ADDR_WIDTH                             : natural;
    BUS_DATA_WIDTH                             : natural;
    BUS_STROBE_WIDTH                           : natural;
    BUS_LEN_WIDTH                              : natural;
    BUS_BURST_STEP_LEN                         : natural;
    BUS_BURST_MAX_LEN                          : natural;
    ---------------------------------------------------------------------------
    INDEX_WIDTH                                : natural;
    ---------------------------------------------------------------------------
    NUM_ARROW_BUFFERS                          : natural;
    NUM_REGS                                   : natural;
    NUM_USER_REGS                              : natural;
    REG_WIDTH                                  : natural;
    ---------------------------------------------------------------------------
    TAG_WIDTH                                  : natural
  );
  port(
    acc_reset                                  : in std_logic;
    bus_clk                                    : in std_logic;
    bus_reset                                  : in std_logic;
    acc_clk                                    : in std_logic;
    ---------------------------------------------------------------------------
    mst_rreq_valid                             : out std_logic;
    mst_rreq_ready                             : in std_logic;
    mst_rreq_addr                              : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    mst_rreq_len                               : out std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
    ---------------------------------------------------------------------------
    mst_rdat_valid                             : in std_logic;
    mst_rdat_ready                             : out std_logic;
    mst_rdat_data                              : in std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
    mst_rdat_last                              : in std_logic;
    ---------------------------------------------------------------------------
    mst_wreq_valid                             : out std_logic;
    mst_wreq_len                               : out std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
    mst_wreq_addr                              : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    mst_wreq_ready                             : in std_logic;
    ---------------------------------------------------------------------------
    mst_wdat_valid                             : out std_logic;
    mst_wdat_ready                             : in std_logic;
    mst_wdat_data                              : out std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
    mst_wdat_strobe                            : out std_logic_vector(BUS_STROBE_WIDTH-1 downto 0);
    mst_wdat_last                              : out std_logic;
    ---------------------------------------------------------------------------
    regs_in                                    : in std_logic_vector(NUM_REGS*REG_WIDTH-1 downto 0);
    regs_out                                   : out std_logic_vector(NUM_REGS*REG_WIDTH-1 downto 0);
    regs_out_en                                : out std_logic_vector(NUM_REGS-1 downto 0)
  );
end fletcher_wrapper;

architecture Implementation of fletcher_wrapper is

  -----------------------------------------------------------------------------
  -- Hardware Accelerated Function component.
  -- This component should be implemented by the user.
  component sum is
    generic(
      TAG_WIDTH                                  : natural;
      BUS_ADDR_WIDTH                             : natural;
      INDEX_WIDTH                                : natural;
      REG_WIDTH                                  : natural
    );
    port(
      weight4_out_last                           : in std_logic;
      weight5_out_last                           : in std_logic;
      weight5_out_ready                          : out std_logic;
      weight5_out_valid                          : in std_logic;
      weight4_cmd_weight4_values_addr            : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      weight4_cmd_tag                            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      weight4_cmd_lastIdx                        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      weight4_cmd_firstIdx                       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      weight4_cmd_ready                          : in std_logic;
      weight4_cmd_valid                          : out std_logic;
      weight4_out_data                           : in std_logic_vector(63 downto 0);
      weight5_out_data                           : in std_logic_vector(63 downto 0);
      weight4_out_ready                          : out std_logic;
      weight4_out_valid                          : in std_logic;
      weight3_cmd_weight3_values_addr            : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      weight3_cmd_tag                            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      weight3_cmd_lastIdx                        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      weight3_cmd_firstIdx                       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      weight3_cmd_ready                          : in std_logic;
      weight3_cmd_valid                          : out std_logic;
      weight3_out_data                           : in std_logic_vector(63 downto 0);
      weight6_out_data                           : in std_logic_vector(63 downto 0);
      weight7_out_last                           : in std_logic;
      weight7_out_ready                          : out std_logic;
      weight7_out_valid                          : in std_logic;
      weight6_cmd_weight6_values_addr            : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      weight6_cmd_tag                            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      weight6_cmd_lastIdx                        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      weight6_cmd_firstIdx                       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      weight6_cmd_ready                          : in std_logic;
      weight6_cmd_valid                          : out std_logic;
      weight3_out_last                           : in std_logic;
      weight6_out_last                           : in std_logic;
      weight6_out_ready                          : out std_logic;
      weight6_out_valid                          : in std_logic;
      weight5_cmd_weight5_values_addr            : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      weight5_cmd_tag                            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      weight5_cmd_lastIdx                        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      weight5_cmd_firstIdx                       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      weight5_cmd_ready                          : in std_logic;
      weight5_cmd_valid                          : out std_logic;
      weight0_out_last                           : in std_logic;
      weight1_out_ready                          : out std_logic;
      weight1_out_valid                          : in std_logic;
      weight0_cmd_weight0_values_addr            : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      weight0_cmd_tag                            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      weight0_cmd_lastIdx                        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      weight0_cmd_firstIdx                       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      weight0_cmd_ready                          : in std_logic;
      weight0_cmd_valid                          : out std_logic;
      weight0_out_data                           : in std_logic_vector(63 downto 0);
      weight1_out_last                           : in std_logic;
      weight0_out_ready                          : out std_logic;
      weight0_out_valid                          : in std_logic;
      weight7_out_data                           : in std_logic_vector(63 downto 0);
      weight7_cmd_valid                          : out std_logic;
      weight7_cmd_ready                          : in std_logic;
      weight7_cmd_firstIdx                       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      weight7_cmd_lastIdx                        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      weight7_cmd_tag                            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      weight7_cmd_weight7_values_addr            : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      weight2_out_last                           : in std_logic;
      weight3_out_ready                          : out std_logic;
      weight3_out_valid                          : in std_logic;
      weight2_cmd_weight2_values_addr            : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      weight2_cmd_tag                            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      weight2_cmd_lastIdx                        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      weight2_cmd_firstIdx                       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      weight2_cmd_ready                          : in std_logic;
      weight2_cmd_valid                          : out std_logic;
      weight2_out_data                           : in std_logic_vector(63 downto 0);
      weight2_out_ready                          : out std_logic;
      weight2_out_valid                          : in std_logic;
      weight1_cmd_weight1_values_addr            : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      weight1_cmd_tag                            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      weight1_cmd_lastIdx                        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      weight1_cmd_firstIdx                       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      weight1_cmd_ready                          : in std_logic;
      weight1_cmd_valid                          : out std_logic;
      weight1_out_data                           : in std_logic_vector(63 downto 0);
      -------------------------------------------------------------------------
      acc_reset                                  : in std_logic;
      acc_clk                                    : in std_logic;
      -------------------------------------------------------------------------
      ctrl_busy                                  : out std_logic;
      ctrl_idle                                  : out std_logic;
      ctrl_reset                                 : in std_logic;
      ctrl_stop                                  : in std_logic;
      ctrl_start                                 : in std_logic;
      ctrl_done                                  : out std_logic;
      -------------------------------------------------------------------------
      reg_return0                                : out std_logic_vector(REG_WIDTH-1 downto 0);
      reg_return1                                : out std_logic_vector(REG_WIDTH-1 downto 0);
      idx_last                                   : in std_logic_vector(REG_WIDTH-1 downto 0);
      idx_first                                  : in std_logic_vector(REG_WIDTH-1 downto 0);
      -------------------------------------------------------------------------
      reg_weight0_values_addr                    : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      reg_weight1_values_addr                    : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      reg_weight2_values_addr                    : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      reg_weight3_values_addr                    : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      reg_weight4_values_addr                    : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      reg_weight5_values_addr                    : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      reg_weight6_values_addr                    : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      reg_weight7_values_addr                    : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0)
    );
  end component;
  -----------------------------------------------------------------------------

  signal s_weight0_cmd_ready                   : std_logic;
  signal uctrl_done                            : std_logic;
  signal uctrl_busy                            : std_logic;
  signal uctrl_idle                            : std_logic;
  signal uctrl_reset                           : std_logic;
  signal uctrl_stop                            : std_logic;
  signal uctrl_start                           : std_logic;
  signal uctrl_control                         : std_logic_vector(REG_WIDTH-1 downto 0);
  signal uctrl_status                          : std_logic_vector(REG_WIDTH-1 downto 0);
  signal s_weight0_bus_rdat_last               : std_logic;
  signal s_weight0_bus_rdat_data               : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal s_weight0_bus_rdat_ready              : std_logic;
  signal s_weight0_bus_rdat_valid              : std_logic;
  signal s_weight0_bus_rreq_len                : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal s_weight0_bus_rreq_ready              : std_logic;
  signal s_weight0_cmd_valid                   : std_logic;
  signal s_weight0_cmd_firstIdx                : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_weight0_cmd_lastIdx                 : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_weight0_cmd_ctrl                    : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_weight0_cmd_tag                     : std_logic_vector(TAG_WIDTH-1 downto 0);
  signal s_weight0_out_valid                   : std_logic_vector(0 downto 0);
  signal s_weight0_out_ready                   : std_logic_vector(0 downto 0);
  signal s_weight0_out_last                    : std_logic_vector(0 downto 0);
  signal s_weight0_bus_rreq_addr               : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_weight0_bus_rreq_valid              : std_logic;
  signal s_weight0_out_dvalid                  : std_logic_vector(0 downto 0);
  signal s_weight0_out_data                    : std_logic_vector(63 downto 0);
  -----------------------------------------------------------------------------
  signal s_weight1_cmd_tag                     : std_logic_vector(TAG_WIDTH-1 downto 0);
  signal s_weight1_cmd_valid                   : std_logic;
  signal s_weight1_cmd_ready                   : std_logic;
  signal s_weight1_cmd_firstIdx                : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_weight1_cmd_lastIdx                 : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_weight1_bus_rdat_last               : std_logic;
  signal s_weight1_bus_rdat_data               : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal s_weight1_bus_rdat_ready              : std_logic;
  signal s_weight1_bus_rreq_len                : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal s_weight1_cmd_ctrl                    : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_weight1_out_valid                   : std_logic_vector(0 downto 0);
  signal s_weight1_out_ready                   : std_logic_vector(0 downto 0);
  signal s_weight1_out_last                    : std_logic_vector(0 downto 0);
  signal s_weight1_out_data                    : std_logic_vector(63 downto 0);
  signal s_weight1_out_dvalid                  : std_logic_vector(0 downto 0);
  signal s_weight1_bus_rreq_valid              : std_logic;
  signal s_weight1_bus_rreq_ready              : std_logic;
  signal s_weight1_bus_rdat_valid              : std_logic;
  signal s_weight1_bus_rreq_addr               : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  -----------------------------------------------------------------------------
  signal s_weight2_out_ready                   : std_logic_vector(0 downto 0);
  signal s_weight2_cmd_valid                   : std_logic;
  signal s_weight2_cmd_ready                   : std_logic;
  signal s_weight2_cmd_firstIdx                : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_weight2_cmd_lastIdx                 : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_weight2_cmd_ctrl                    : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_weight2_cmd_tag                     : std_logic_vector(TAG_WIDTH-1 downto 0);
  signal s_weight2_bus_rdat_last               : std_logic;
  signal s_weight2_bus_rdat_data               : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal s_weight2_bus_rdat_valid              : std_logic;
  signal s_weight2_out_valid                   : std_logic_vector(0 downto 0);
  signal s_weight2_out_last                    : std_logic_vector(0 downto 0);
  signal s_weight2_out_data                    : std_logic_vector(63 downto 0);
  signal s_weight2_out_dvalid                  : std_logic_vector(0 downto 0);
  signal s_weight2_bus_rreq_valid              : std_logic;
  signal s_weight2_bus_rreq_ready              : std_logic;
  signal s_weight2_bus_rreq_addr               : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_weight2_bus_rreq_len                : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal s_weight2_bus_rdat_ready              : std_logic;
  -----------------------------------------------------------------------------
  signal s_weight3_out_last                    : std_logic_vector(0 downto 0);
  signal s_weight3_cmd_valid                   : std_logic;
  signal s_weight3_cmd_ready                   : std_logic;
  signal s_weight3_cmd_firstIdx                : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_weight3_cmd_lastIdx                 : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_weight3_cmd_ctrl                    : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_weight3_cmd_tag                     : std_logic_vector(TAG_WIDTH-1 downto 0);
  signal s_weight3_out_valid                   : std_logic_vector(0 downto 0);
  signal s_weight3_bus_rdat_last               : std_logic;
  signal s_weight3_bus_rdat_ready              : std_logic;
  signal s_weight3_out_ready                   : std_logic_vector(0 downto 0);
  signal s_weight3_out_data                    : std_logic_vector(63 downto 0);
  signal s_weight3_out_dvalid                  : std_logic_vector(0 downto 0);
  signal s_weight3_bus_rreq_valid              : std_logic;
  signal s_weight3_bus_rreq_ready              : std_logic;
  signal s_weight3_bus_rreq_addr               : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_weight3_bus_rreq_len                : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal s_weight3_bus_rdat_valid              : std_logic;
  signal s_weight3_bus_rdat_data               : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  -----------------------------------------------------------------------------
  signal s_weight4_out_last                    : std_logic_vector(0 downto 0);
  signal s_weight4_cmd_valid                   : std_logic;
  signal s_weight4_cmd_ready                   : std_logic;
  signal s_weight4_cmd_firstIdx                : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_weight4_cmd_lastIdx                 : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_weight4_cmd_ctrl                    : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_weight4_cmd_tag                     : std_logic_vector(TAG_WIDTH-1 downto 0);
  signal s_weight4_out_valid                   : std_logic_vector(0 downto 0);
  signal s_weight4_bus_rdat_last               : std_logic;
  signal s_weight4_bus_rdat_ready              : std_logic;
  signal s_weight4_out_ready                   : std_logic_vector(0 downto 0);
  signal s_weight4_out_data                    : std_logic_vector(63 downto 0);
  signal s_weight4_out_dvalid                  : std_logic_vector(0 downto 0);
  signal s_weight4_bus_rreq_valid              : std_logic;
  signal s_weight4_bus_rreq_ready              : std_logic;
  signal s_weight4_bus_rreq_addr               : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_weight4_bus_rreq_len                : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal s_weight4_bus_rdat_valid              : std_logic;
  signal s_weight4_bus_rdat_data               : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  -----------------------------------------------------------------------------
  signal s_weight5_out_last                    : std_logic_vector(0 downto 0);
  signal s_weight5_cmd_valid                   : std_logic;
  signal s_weight5_cmd_ready                   : std_logic;
  signal s_weight5_cmd_firstIdx                : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_weight5_cmd_lastIdx                 : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_weight5_cmd_ctrl                    : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_weight5_cmd_tag                     : std_logic_vector(TAG_WIDTH-1 downto 0);
  signal s_weight5_out_valid                   : std_logic_vector(0 downto 0);
  signal s_weight5_bus_rdat_last               : std_logic;
  signal s_weight5_bus_rdat_ready              : std_logic;
  signal s_weight5_out_ready                   : std_logic_vector(0 downto 0);
  signal s_weight5_out_data                    : std_logic_vector(63 downto 0);
  signal s_weight5_out_dvalid                  : std_logic_vector(0 downto 0);
  signal s_weight5_bus_rreq_valid              : std_logic;
  signal s_weight5_bus_rreq_ready              : std_logic;
  signal s_weight5_bus_rreq_addr               : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_weight5_bus_rreq_len                : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal s_weight5_bus_rdat_valid              : std_logic;
  signal s_weight5_bus_rdat_data               : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  -----------------------------------------------------------------------------
  signal s_weight6_out_last                    : std_logic_vector(0 downto 0);
  signal s_weight6_cmd_valid                   : std_logic;
  signal s_weight6_cmd_ready                   : std_logic;
  signal s_weight6_cmd_firstIdx                : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_weight6_cmd_lastIdx                 : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_weight6_cmd_ctrl                    : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_weight6_cmd_tag                     : std_logic_vector(TAG_WIDTH-1 downto 0);
  signal s_weight6_out_valid                   : std_logic_vector(0 downto 0);
  signal s_weight6_bus_rdat_last               : std_logic;
  signal s_weight6_bus_rdat_ready              : std_logic;
  signal s_weight6_out_ready                   : std_logic_vector(0 downto 0);
  signal s_weight6_out_data                    : std_logic_vector(63 downto 0);
  signal s_weight6_out_dvalid                  : std_logic_vector(0 downto 0);
  signal s_weight6_bus_rreq_valid              : std_logic;
  signal s_weight6_bus_rreq_ready              : std_logic;
  signal s_weight6_bus_rreq_addr               : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_weight6_bus_rreq_len                : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal s_weight6_bus_rdat_valid              : std_logic;
  signal s_weight6_bus_rdat_data               : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  -----------------------------------------------------------------------------
  signal s_weight7_bus_rdat_data               : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal s_weight7_bus_rdat_valid              : std_logic;
  signal s_weight7_cmd_ctrl                    : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_weight7_bus_rreq_len                : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal s_weight7_out_ready                   : std_logic_vector(0 downto 0);
  signal s_weight7_out_valid                   : std_logic_vector(0 downto 0);
  signal s_weight7_cmd_tag                     : std_logic_vector(TAG_WIDTH-1 downto 0);
  signal s_weight7_cmd_lastIdx                 : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_weight7_cmd_firstIdx                : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_weight7_cmd_valid                   : std_logic;
  signal s_weight7_out_data                    : std_logic_vector(63 downto 0);
  signal s_weight7_bus_rreq_ready              : std_logic;
  signal s_weight7_out_dvalid                  : std_logic_vector(0 downto 0);
  signal s_weight7_cmd_ready                   : std_logic;
  signal s_weight7_bus_rdat_ready              : std_logic;
  signal s_weight7_bus_rreq_valid              : std_logic;
  signal s_weight7_out_last                    : std_logic_vector(0 downto 0);
  signal s_weight7_bus_rdat_last               : std_logic;
  signal s_weight7_bus_rreq_addr               : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  -----------------------------------------------------------------------------
  signal s_bsv_rreq_len                        : std_logic_vector(8*BUS_LEN_WIDTH-1 downto 0);
  signal s_bsv_rreq_valid                      : std_logic_vector(7 downto 0);
  signal s_bsv_rreq_ready                      : std_logic_vector(7 downto 0);
  signal s_bsv_rreq_addr                       : std_logic_vector(8*BUS_ADDR_WIDTH-1 downto 0);
  -----------------------------------------------------------------------------
  signal s_bsv_rdat_valid                      : std_logic_vector(7 downto 0);
  signal s_bsv_rdat_ready                      : std_logic_vector(7 downto 0);
  signal s_bsv_rdat_data                       : std_logic_vector(8*BUS_DATA_WIDTH-1 downto 0);
  signal s_bsv_rdat_last                       : std_logic_vector(7 downto 0);
begin
  -- ColumnReader instance generated from Arrow schema field:
  -- weight0: int64 not null
  weight0_read_inst: ColumnReader
    generic map (
      CFG                                      => "prim(64)",
      BUS_ADDR_WIDTH                           => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH                            => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH                           => BUS_DATA_WIDTH,
      BUS_BURST_STEP_LEN                       => BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN                        => BUS_BURST_MAX_LEN,
      INDEX_WIDTH                              => INDEX_WIDTH
    )
    port map (
      bus_clk                                  => bus_clk,
      bus_reset                                => bus_reset,
      acc_clk                                  => acc_clk,
      acc_reset                                => acc_reset,
      cmd_valid                                => s_weight0_cmd_valid,
      cmd_ready                                => s_weight0_cmd_ready,
      cmd_firstIdx                             => s_weight0_cmd_firstIdx,
      cmd_lastIdx                              => s_weight0_cmd_lastIdx,
      cmd_ctrl                                 => s_weight0_cmd_ctrl,
      cmd_tag                                  => s_weight0_cmd_tag,
      out_valid                                => s_weight0_out_valid,
      out_ready                                => s_weight0_out_ready,
      out_last                                 => s_weight0_out_last,
      out_data                                 => s_weight0_out_data,
      out_dvalid                               => s_weight0_out_dvalid,
      bus_rreq_valid                           => s_weight0_bus_rreq_valid,
      bus_rreq_ready                           => s_weight0_bus_rreq_ready,
      bus_rreq_addr                            => s_weight0_bus_rreq_addr,
      bus_rreq_len                             => s_weight0_bus_rreq_len,
      bus_rdat_valid                           => s_weight0_bus_rdat_valid,
      bus_rdat_ready                           => s_weight0_bus_rdat_ready,
      bus_rdat_data                            => s_weight0_bus_rdat_data,
      bus_rdat_last                            => s_weight0_bus_rdat_last
    );

  -- ColumnReader instance generated from Arrow schema field:
  -- weight1: int64 not null
  weight1_read_inst: ColumnReader
    generic map (
      CFG                                      => "prim(64)",
      BUS_ADDR_WIDTH                           => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH                            => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH                           => BUS_DATA_WIDTH,
      BUS_BURST_STEP_LEN                       => BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN                        => BUS_BURST_MAX_LEN,
      INDEX_WIDTH                              => INDEX_WIDTH
    )
    port map (
      bus_clk                                  => bus_clk,
      bus_reset                                => bus_reset,
      acc_clk                                  => acc_clk,
      acc_reset                                => acc_reset,
      cmd_valid                                => s_weight1_cmd_valid,
      cmd_ready                                => s_weight1_cmd_ready,
      cmd_firstIdx                             => s_weight1_cmd_firstIdx,
      cmd_lastIdx                              => s_weight1_cmd_lastIdx,
      cmd_ctrl                                 => s_weight1_cmd_ctrl,
      cmd_tag                                  => s_weight1_cmd_tag,
      out_valid                                => s_weight1_out_valid,
      out_ready                                => s_weight1_out_ready,
      out_last                                 => s_weight1_out_last,
      out_data                                 => s_weight1_out_data,
      out_dvalid                               => s_weight1_out_dvalid,
      bus_rreq_valid                           => s_weight1_bus_rreq_valid,
      bus_rreq_ready                           => s_weight1_bus_rreq_ready,
      bus_rreq_addr                            => s_weight1_bus_rreq_addr,
      bus_rreq_len                             => s_weight1_bus_rreq_len,
      bus_rdat_valid                           => s_weight1_bus_rdat_valid,
      bus_rdat_ready                           => s_weight1_bus_rdat_ready,
      bus_rdat_data                            => s_weight1_bus_rdat_data,
      bus_rdat_last                            => s_weight1_bus_rdat_last
    );

  -- ColumnReader instance generated from Arrow schema field:
  -- weight2: int64 not null
  weight2_read_inst: ColumnReader
    generic map (
      CFG                                      => "prim(64)",
      BUS_ADDR_WIDTH                           => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH                            => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH                           => BUS_DATA_WIDTH,
      BUS_BURST_STEP_LEN                       => BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN                        => BUS_BURST_MAX_LEN,
      INDEX_WIDTH                              => INDEX_WIDTH
    )
    port map (
      bus_clk                                  => bus_clk,
      bus_reset                                => bus_reset,
      acc_clk                                  => acc_clk,
      acc_reset                                => acc_reset,
      cmd_valid                                => s_weight2_cmd_valid,
      cmd_ready                                => s_weight2_cmd_ready,
      cmd_firstIdx                             => s_weight2_cmd_firstIdx,
      cmd_lastIdx                              => s_weight2_cmd_lastIdx,
      cmd_ctrl                                 => s_weight2_cmd_ctrl,
      cmd_tag                                  => s_weight2_cmd_tag,
      out_valid                                => s_weight2_out_valid,
      out_ready                                => s_weight2_out_ready,
      out_last                                 => s_weight2_out_last,
      out_data                                 => s_weight2_out_data,
      out_dvalid                               => s_weight2_out_dvalid,
      bus_rreq_valid                           => s_weight2_bus_rreq_valid,
      bus_rreq_ready                           => s_weight2_bus_rreq_ready,
      bus_rreq_addr                            => s_weight2_bus_rreq_addr,
      bus_rreq_len                             => s_weight2_bus_rreq_len,
      bus_rdat_valid                           => s_weight2_bus_rdat_valid,
      bus_rdat_ready                           => s_weight2_bus_rdat_ready,
      bus_rdat_data                            => s_weight2_bus_rdat_data,
      bus_rdat_last                            => s_weight2_bus_rdat_last
    );

  -- ColumnReader instance generated from Arrow schema field:
  -- weight3: int64 not null
  weight3_read_inst: ColumnReader
    generic map (
      CFG                                      => "prim(64)",
      BUS_ADDR_WIDTH                           => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH                            => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH                           => BUS_DATA_WIDTH,
      BUS_BURST_STEP_LEN                       => BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN                        => BUS_BURST_MAX_LEN,
      INDEX_WIDTH                              => INDEX_WIDTH
    )
    port map (
      bus_clk                                  => bus_clk,
      bus_reset                                => bus_reset,
      acc_clk                                  => acc_clk,
      acc_reset                                => acc_reset,
      cmd_valid                                => s_weight3_cmd_valid,
      cmd_ready                                => s_weight3_cmd_ready,
      cmd_firstIdx                             => s_weight3_cmd_firstIdx,
      cmd_lastIdx                              => s_weight3_cmd_lastIdx,
      cmd_ctrl                                 => s_weight3_cmd_ctrl,
      cmd_tag                                  => s_weight3_cmd_tag,
      out_valid                                => s_weight3_out_valid,
      out_ready                                => s_weight3_out_ready,
      out_last                                 => s_weight3_out_last,
      out_data                                 => s_weight3_out_data,
      out_dvalid                               => s_weight3_out_dvalid,
      bus_rreq_valid                           => s_weight3_bus_rreq_valid,
      bus_rreq_ready                           => s_weight3_bus_rreq_ready,
      bus_rreq_addr                            => s_weight3_bus_rreq_addr,
      bus_rreq_len                             => s_weight3_bus_rreq_len,
      bus_rdat_valid                           => s_weight3_bus_rdat_valid,
      bus_rdat_ready                           => s_weight3_bus_rdat_ready,
      bus_rdat_data                            => s_weight3_bus_rdat_data,
      bus_rdat_last                            => s_weight3_bus_rdat_last
    );

  -- ColumnReader instance generated from Arrow schema field:
  -- weight4: int64 not null
  weight4_read_inst: ColumnReader
    generic map (
      CFG                                      => "prim(64)",
      BUS_ADDR_WIDTH                           => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH                            => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH                           => BUS_DATA_WIDTH,
      BUS_BURST_STEP_LEN                       => BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN                        => BUS_BURST_MAX_LEN,
      INDEX_WIDTH                              => INDEX_WIDTH
    )
    port map (
      bus_clk                                  => bus_clk,
      bus_reset                                => bus_reset,
      acc_clk                                  => acc_clk,
      acc_reset                                => acc_reset,
      cmd_valid                                => s_weight4_cmd_valid,
      cmd_ready                                => s_weight4_cmd_ready,
      cmd_firstIdx                             => s_weight4_cmd_firstIdx,
      cmd_lastIdx                              => s_weight4_cmd_lastIdx,
      cmd_ctrl                                 => s_weight4_cmd_ctrl,
      cmd_tag                                  => s_weight4_cmd_tag,
      out_valid                                => s_weight4_out_valid,
      out_ready                                => s_weight4_out_ready,
      out_last                                 => s_weight4_out_last,
      out_data                                 => s_weight4_out_data,
      out_dvalid                               => s_weight4_out_dvalid,
      bus_rreq_valid                           => s_weight4_bus_rreq_valid,
      bus_rreq_ready                           => s_weight4_bus_rreq_ready,
      bus_rreq_addr                            => s_weight4_bus_rreq_addr,
      bus_rreq_len                             => s_weight4_bus_rreq_len,
      bus_rdat_valid                           => s_weight4_bus_rdat_valid,
      bus_rdat_ready                           => s_weight4_bus_rdat_ready,
      bus_rdat_data                            => s_weight4_bus_rdat_data,
      bus_rdat_last                            => s_weight4_bus_rdat_last
    );

  -- ColumnReader instance generated from Arrow schema field:
  -- weight5: int64 not null
  weight5_read_inst: ColumnReader
    generic map (
      CFG                                      => "prim(64)",
      BUS_ADDR_WIDTH                           => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH                            => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH                           => BUS_DATA_WIDTH,
      BUS_BURST_STEP_LEN                       => BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN                        => BUS_BURST_MAX_LEN,
      INDEX_WIDTH                              => INDEX_WIDTH
    )
    port map (
      bus_clk                                  => bus_clk,
      bus_reset                                => bus_reset,
      acc_clk                                  => acc_clk,
      acc_reset                                => acc_reset,
      cmd_valid                                => s_weight5_cmd_valid,
      cmd_ready                                => s_weight5_cmd_ready,
      cmd_firstIdx                             => s_weight5_cmd_firstIdx,
      cmd_lastIdx                              => s_weight5_cmd_lastIdx,
      cmd_ctrl                                 => s_weight5_cmd_ctrl,
      cmd_tag                                  => s_weight5_cmd_tag,
      out_valid                                => s_weight5_out_valid,
      out_ready                                => s_weight5_out_ready,
      out_last                                 => s_weight5_out_last,
      out_data                                 => s_weight5_out_data,
      out_dvalid                               => s_weight5_out_dvalid,
      bus_rreq_valid                           => s_weight5_bus_rreq_valid,
      bus_rreq_ready                           => s_weight5_bus_rreq_ready,
      bus_rreq_addr                            => s_weight5_bus_rreq_addr,
      bus_rreq_len                             => s_weight5_bus_rreq_len,
      bus_rdat_valid                           => s_weight5_bus_rdat_valid,
      bus_rdat_ready                           => s_weight5_bus_rdat_ready,
      bus_rdat_data                            => s_weight5_bus_rdat_data,
      bus_rdat_last                            => s_weight5_bus_rdat_last
    );

  -- ColumnReader instance generated from Arrow schema field:
  -- weight6: int64 not null
  weight6_read_inst: ColumnReader
    generic map (
      CFG                                      => "prim(64)",
      BUS_ADDR_WIDTH                           => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH                            => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH                           => BUS_DATA_WIDTH,
      BUS_BURST_STEP_LEN                       => BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN                        => BUS_BURST_MAX_LEN,
      INDEX_WIDTH                              => INDEX_WIDTH
    )
    port map (
      bus_clk                                  => bus_clk,
      bus_reset                                => bus_reset,
      acc_clk                                  => acc_clk,
      acc_reset                                => acc_reset,
      cmd_valid                                => s_weight6_cmd_valid,
      cmd_ready                                => s_weight6_cmd_ready,
      cmd_firstIdx                             => s_weight6_cmd_firstIdx,
      cmd_lastIdx                              => s_weight6_cmd_lastIdx,
      cmd_ctrl                                 => s_weight6_cmd_ctrl,
      cmd_tag                                  => s_weight6_cmd_tag,
      out_valid                                => s_weight6_out_valid,
      out_ready                                => s_weight6_out_ready,
      out_last                                 => s_weight6_out_last,
      out_data                                 => s_weight6_out_data,
      out_dvalid                               => s_weight6_out_dvalid,
      bus_rreq_valid                           => s_weight6_bus_rreq_valid,
      bus_rreq_ready                           => s_weight6_bus_rreq_ready,
      bus_rreq_addr                            => s_weight6_bus_rreq_addr,
      bus_rreq_len                             => s_weight6_bus_rreq_len,
      bus_rdat_valid                           => s_weight6_bus_rdat_valid,
      bus_rdat_ready                           => s_weight6_bus_rdat_ready,
      bus_rdat_data                            => s_weight6_bus_rdat_data,
      bus_rdat_last                            => s_weight6_bus_rdat_last
    );

  -- ColumnReader instance generated from Arrow schema field:
  -- weight7: int64 not null
  weight7_read_inst: ColumnReader
    generic map (
      CFG                                      => "prim(64)",
      BUS_ADDR_WIDTH                           => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH                            => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH                           => BUS_DATA_WIDTH,
      BUS_BURST_STEP_LEN                       => BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN                        => BUS_BURST_MAX_LEN,
      INDEX_WIDTH                              => INDEX_WIDTH
    )
    port map (
      bus_clk                                  => bus_clk,
      bus_reset                                => bus_reset,
      acc_clk                                  => acc_clk,
      acc_reset                                => acc_reset,
      cmd_valid                                => s_weight7_cmd_valid,
      cmd_ready                                => s_weight7_cmd_ready,
      cmd_firstIdx                             => s_weight7_cmd_firstIdx,
      cmd_lastIdx                              => s_weight7_cmd_lastIdx,
      cmd_ctrl                                 => s_weight7_cmd_ctrl,
      cmd_tag                                  => s_weight7_cmd_tag,
      out_valid                                => s_weight7_out_valid,
      out_ready                                => s_weight7_out_ready,
      out_last                                 => s_weight7_out_last,
      out_data                                 => s_weight7_out_data,
      out_dvalid                               => s_weight7_out_dvalid,
      bus_rreq_valid                           => s_weight7_bus_rreq_valid,
      bus_rreq_ready                           => s_weight7_bus_rreq_ready,
      bus_rreq_addr                            => s_weight7_bus_rreq_addr,
      bus_rreq_len                             => s_weight7_bus_rreq_len,
      bus_rdat_valid                           => s_weight7_bus_rdat_valid,
      bus_rdat_ready                           => s_weight7_bus_rdat_ready,
      bus_rdat_data                            => s_weight7_bus_rdat_data,
      bus_rdat_last                            => s_weight7_bus_rdat_last
    );

  -- Controller instance.
  UserCoreController_inst: UserCoreController
    generic map (
      REG_WIDTH                                => REG_WIDTH
    )
    port map (
      acc_clk                                  => acc_clk,
      acc_reset                                => acc_reset,
      bus_clk                                  => bus_clk,
      bus_reset                                => bus_reset,
      status                                   => regs_out(2*REG_WIDTH-1 downto REG_WIDTH),
      control                                  => regs_in(REG_WIDTH-1 downto 0),
      start                                    => uctrl_start,
      stop                                     => uctrl_stop,
      reset                                    => uctrl_reset,
      idle                                     => uctrl_idle,
      busy                                     => uctrl_busy,
      done                                     => uctrl_done
    );

  -- Hardware Accelerated Function instance.
  sum_inst: sum
    generic map (
      TAG_WIDTH                                => TAG_WIDTH,
      BUS_ADDR_WIDTH                           => BUS_ADDR_WIDTH,
      INDEX_WIDTH                              => INDEX_WIDTH,
      REG_WIDTH                                => REG_WIDTH
    )
    port map (
      acc_clk                                  => acc_clk,
      acc_reset                                => acc_reset,
      ctrl_start                               => uctrl_start,
      ctrl_stop                                => uctrl_stop,
      ctrl_reset                               => uctrl_reset,
      ctrl_idle                                => uctrl_idle,
      ctrl_busy                                => uctrl_busy,
      ctrl_done                                => uctrl_done,
      weight0_out_valid                        => s_weight0_out_valid(0),
      weight0_out_ready                        => s_weight0_out_ready(0),
      weight0_out_last                         => s_weight0_out_last(0),
      weight0_out_data                         => s_weight0_out_data(63 downto 0),
      weight0_cmd_valid                        => s_weight0_cmd_valid,
      weight0_cmd_ready                        => s_weight0_cmd_ready,
      weight0_cmd_firstIdx                     => s_weight0_cmd_firstIdx(INDEX_WIDTH-1 downto 0),
      weight0_cmd_lastIdx                      => s_weight0_cmd_lastIdx(INDEX_WIDTH-1 downto 0),
      weight0_cmd_tag                          => s_weight0_cmd_tag(TAG_WIDTH-1 downto 0),
      weight0_cmd_weight0_values_addr          => s_weight0_cmd_ctrl(BUS_ADDR_WIDTH-1 downto 0),
      weight1_out_valid                        => s_weight1_out_valid(0),
      weight1_out_ready                        => s_weight1_out_ready(0),
      weight1_out_last                         => s_weight1_out_last(0),
      weight1_out_data                         => s_weight1_out_data(63 downto 0),
      weight1_cmd_valid                        => s_weight1_cmd_valid,
      weight1_cmd_ready                        => s_weight1_cmd_ready,
      weight1_cmd_firstIdx                     => s_weight1_cmd_firstIdx(INDEX_WIDTH-1 downto 0),
      weight1_cmd_lastIdx                      => s_weight1_cmd_lastIdx(INDEX_WIDTH-1 downto 0),
      weight1_cmd_tag                          => s_weight1_cmd_tag(TAG_WIDTH-1 downto 0),
      weight1_cmd_weight1_values_addr          => s_weight1_cmd_ctrl(BUS_ADDR_WIDTH-1 downto 0),
      weight2_out_valid                        => s_weight2_out_valid(0),
      weight2_out_ready                        => s_weight2_out_ready(0),
      weight2_out_last                         => s_weight2_out_last(0),
      weight2_out_data                         => s_weight2_out_data(63 downto 0),
      weight2_cmd_valid                        => s_weight2_cmd_valid,
      weight2_cmd_ready                        => s_weight2_cmd_ready,
      weight2_cmd_firstIdx                     => s_weight2_cmd_firstIdx(INDEX_WIDTH-1 downto 0),
      weight2_cmd_lastIdx                      => s_weight2_cmd_lastIdx(INDEX_WIDTH-1 downto 0),
      weight2_cmd_tag                          => s_weight2_cmd_tag(TAG_WIDTH-1 downto 0),
      weight2_cmd_weight2_values_addr          => s_weight2_cmd_ctrl(BUS_ADDR_WIDTH-1 downto 0),
      weight3_out_valid                        => s_weight3_out_valid(0),
      weight3_out_ready                        => s_weight3_out_ready(0),
      weight3_out_last                         => s_weight3_out_last(0),
      weight3_out_data                         => s_weight3_out_data(63 downto 0),
      weight3_cmd_valid                        => s_weight3_cmd_valid,
      weight3_cmd_ready                        => s_weight3_cmd_ready,
      weight3_cmd_firstIdx                     => s_weight3_cmd_firstIdx(INDEX_WIDTH-1 downto 0),
      weight3_cmd_lastIdx                      => s_weight3_cmd_lastIdx(INDEX_WIDTH-1 downto 0),
      weight3_cmd_tag                          => s_weight3_cmd_tag(TAG_WIDTH-1 downto 0),
      weight3_cmd_weight3_values_addr          => s_weight3_cmd_ctrl(BUS_ADDR_WIDTH-1 downto 0),
      weight4_out_valid                        => s_weight4_out_valid(0),
      weight4_out_ready                        => s_weight4_out_ready(0),
      weight4_out_last                         => s_weight4_out_last(0),
      weight4_out_data                         => s_weight4_out_data(63 downto 0),
      weight4_cmd_valid                        => s_weight4_cmd_valid,
      weight4_cmd_ready                        => s_weight4_cmd_ready,
      weight4_cmd_firstIdx                     => s_weight4_cmd_firstIdx(INDEX_WIDTH-1 downto 0),
      weight4_cmd_lastIdx                      => s_weight4_cmd_lastIdx(INDEX_WIDTH-1 downto 0),
      weight4_cmd_tag                          => s_weight4_cmd_tag(TAG_WIDTH-1 downto 0),
      weight4_cmd_weight4_values_addr          => s_weight4_cmd_ctrl(BUS_ADDR_WIDTH-1 downto 0),
      weight5_out_valid                        => s_weight5_out_valid(0),
      weight5_out_ready                        => s_weight5_out_ready(0),
      weight5_out_last                         => s_weight5_out_last(0),
      weight5_out_data                         => s_weight5_out_data(63 downto 0),
      weight5_cmd_valid                        => s_weight5_cmd_valid,
      weight5_cmd_ready                        => s_weight5_cmd_ready,
      weight5_cmd_firstIdx                     => s_weight5_cmd_firstIdx(INDEX_WIDTH-1 downto 0),
      weight5_cmd_lastIdx                      => s_weight5_cmd_lastIdx(INDEX_WIDTH-1 downto 0),
      weight5_cmd_tag                          => s_weight5_cmd_tag(TAG_WIDTH-1 downto 0),
      weight5_cmd_weight5_values_addr          => s_weight5_cmd_ctrl(BUS_ADDR_WIDTH-1 downto 0),
      weight6_out_valid                        => s_weight6_out_valid(0),
      weight6_out_ready                        => s_weight6_out_ready(0),
      weight6_out_last                         => s_weight6_out_last(0),
      weight6_out_data                         => s_weight6_out_data(63 downto 0),
      weight6_cmd_valid                        => s_weight6_cmd_valid,
      weight6_cmd_ready                        => s_weight6_cmd_ready,
      weight6_cmd_firstIdx                     => s_weight6_cmd_firstIdx(INDEX_WIDTH-1 downto 0),
      weight6_cmd_lastIdx                      => s_weight6_cmd_lastIdx(INDEX_WIDTH-1 downto 0),
      weight6_cmd_tag                          => s_weight6_cmd_tag(TAG_WIDTH-1 downto 0),
      weight6_cmd_weight6_values_addr          => s_weight6_cmd_ctrl(BUS_ADDR_WIDTH-1 downto 0),
      weight7_out_valid                        => s_weight7_out_valid(0),
      weight7_out_ready                        => s_weight7_out_ready(0),
      weight7_out_last                         => s_weight7_out_last(0),
      weight7_out_data                         => s_weight7_out_data(63 downto 0),
      weight7_cmd_valid                        => s_weight7_cmd_valid,
      weight7_cmd_ready                        => s_weight7_cmd_ready,
      weight7_cmd_firstIdx                     => s_weight7_cmd_firstIdx(INDEX_WIDTH-1 downto 0),
      weight7_cmd_lastIdx                      => s_weight7_cmd_lastIdx(INDEX_WIDTH-1 downto 0),
      weight7_cmd_tag                          => s_weight7_cmd_tag(TAG_WIDTH-1 downto 0),
      weight7_cmd_weight7_values_addr          => s_weight7_cmd_ctrl(BUS_ADDR_WIDTH-1 downto 0),
      idx_first                                => regs_in(5*REG_WIDTH-1 downto 4*REG_WIDTH),
      idx_last                                 => regs_in(6*REG_WIDTH-1 downto 5*REG_WIDTH),
      reg_return0                              => regs_out(3*REG_WIDTH-1 downto 2*REG_WIDTH),
      reg_return1                              => regs_out(4*REG_WIDTH-1 downto 3*REG_WIDTH),
      reg_weight0_values_addr                  => regs_in(8*REG_WIDTH-1 downto 6*REG_WIDTH),
      reg_weight1_values_addr                  => regs_in(10*REG_WIDTH-1 downto 8*REG_WIDTH),
      reg_weight2_values_addr                  => regs_in(12*REG_WIDTH-1 downto 10*REG_WIDTH),
      reg_weight3_values_addr                  => regs_in(14*REG_WIDTH-1 downto 12*REG_WIDTH),
      reg_weight4_values_addr                  => regs_in(16*REG_WIDTH-1 downto 14*REG_WIDTH),
      reg_weight5_values_addr                  => regs_in(18*REG_WIDTH-1 downto 16*REG_WIDTH),
      reg_weight6_values_addr                  => regs_in(20*REG_WIDTH-1 downto 18*REG_WIDTH),
      reg_weight7_values_addr                  => regs_in(22*REG_WIDTH-1 downto 20*REG_WIDTH)
    );

  -- Arbiter instance generated to serve 8 column readers.
  BusReadArbiterVec_inst: BusReadArbiterVec
    generic map (
      BUS_ADDR_WIDTH                           => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH                            => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH                           => BUS_DATA_WIDTH,
      NUM_SLAVE_PORTS                          => 8
    )
    port map (
      bus_clk                                  => bus_clk,
      bus_reset                                => bus_reset,
      bsv_rreq_valid                           => s_bsv_rreq_valid,
      bsv_rreq_ready                           => s_bsv_rreq_ready,
      bsv_rreq_addr                            => s_bsv_rreq_addr,
      bsv_rreq_len                             => s_bsv_rreq_len,
      bsv_rdat_valid                           => s_bsv_rdat_valid,
      bsv_rdat_ready                           => s_bsv_rdat_ready,
      bsv_rdat_data                            => s_bsv_rdat_data,
      bsv_rdat_last                            => s_bsv_rdat_last,
      mst_rreq_valid                           => mst_rreq_valid,
      mst_rreq_ready                           => mst_rreq_ready,
      mst_rreq_addr                            => mst_rreq_addr,
      mst_rreq_len                             => mst_rreq_len,
      mst_rdat_valid                           => mst_rdat_valid,
      mst_rdat_ready                           => mst_rdat_ready,
      mst_rdat_data                            => mst_rdat_data,
      mst_rdat_last                            => mst_rdat_last
    );


  s_bsv_rreq_valid(0)                          <= s_weight0_bus_rreq_valid;
  s_weight0_bus_rreq_ready                     <= s_bsv_rreq_ready(0);
  s_bsv_rreq_len(BUS_LEN_WIDTH-1 downto 0)     <= s_weight0_bus_rreq_len;
  s_bsv_rreq_addr(BUS_ADDR_WIDTH-1 downto 0)   <= s_weight0_bus_rreq_addr;
  -----------------------------------------------------------------------------
  s_bsv_rreq_valid(1)                          <= s_weight1_bus_rreq_valid;
  s_weight1_bus_rreq_ready                     <= s_bsv_rreq_ready(1);
  s_bsv_rreq_len(2*BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH)<= s_weight1_bus_rreq_len;
  s_bsv_rreq_addr(2*BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH)<= s_weight1_bus_rreq_addr;
  -----------------------------------------------------------------------------
  s_bsv_rreq_valid(2)                          <= s_weight2_bus_rreq_valid;
  s_weight2_bus_rreq_ready                     <= s_bsv_rreq_ready(2);
  s_bsv_rreq_len(3*BUS_LEN_WIDTH-1 downto 2*BUS_LEN_WIDTH)<= s_weight2_bus_rreq_len;
  s_bsv_rreq_addr(3*BUS_ADDR_WIDTH-1 downto 2*BUS_ADDR_WIDTH)<= s_weight2_bus_rreq_addr;
  -----------------------------------------------------------------------------
  s_bsv_rreq_addr(4*BUS_ADDR_WIDTH-1 downto 3*BUS_ADDR_WIDTH)<= s_weight3_bus_rreq_addr;
  s_bsv_rreq_valid(3)                          <= s_weight3_bus_rreq_valid;
  s_weight3_bus_rreq_ready                     <= s_bsv_rreq_ready(3);
  s_bsv_rreq_len(4*BUS_LEN_WIDTH-1 downto 3*BUS_LEN_WIDTH)<= s_weight3_bus_rreq_len;
  -----------------------------------------------------------------------------
  s_bsv_rreq_addr(5*BUS_ADDR_WIDTH-1 downto 4*BUS_ADDR_WIDTH)<= s_weight4_bus_rreq_addr;
  s_bsv_rreq_valid(4)                          <= s_weight4_bus_rreq_valid;
  s_bsv_rreq_len(5*BUS_LEN_WIDTH-1 downto 4*BUS_LEN_WIDTH)<= s_weight4_bus_rreq_len;
  s_weight4_bus_rreq_ready                     <= s_bsv_rreq_ready(4);
  -----------------------------------------------------------------------------
  s_bsv_rreq_addr(6*BUS_ADDR_WIDTH-1 downto 5*BUS_ADDR_WIDTH)<= s_weight5_bus_rreq_addr;
  s_bsv_rreq_len(6*BUS_LEN_WIDTH-1 downto 5*BUS_LEN_WIDTH)<= s_weight5_bus_rreq_len;
  s_bsv_rreq_valid(5)                          <= s_weight5_bus_rreq_valid;
  s_weight5_bus_rreq_ready                     <= s_bsv_rreq_ready(5);
  -----------------------------------------------------------------------------
  s_bsv_rreq_addr(7*BUS_ADDR_WIDTH-1 downto 6*BUS_ADDR_WIDTH)<= s_weight6_bus_rreq_addr;
  s_bsv_rreq_len(7*BUS_LEN_WIDTH-1 downto 6*BUS_LEN_WIDTH)<= s_weight6_bus_rreq_len;
  s_weight6_bus_rreq_ready                     <= s_bsv_rreq_ready(6);
  s_bsv_rreq_valid(6)                          <= s_weight6_bus_rreq_valid;
  -----------------------------------------------------------------------------
  s_bsv_rreq_len(8*BUS_LEN_WIDTH-1 downto 7*BUS_LEN_WIDTH)<= s_weight7_bus_rreq_len;
  s_weight7_bus_rreq_ready                     <= s_bsv_rreq_ready(7);
  s_bsv_rreq_valid(7)                          <= s_weight7_bus_rreq_valid;
  s_bsv_rreq_addr(8*BUS_ADDR_WIDTH-1 downto 7*BUS_ADDR_WIDTH)<= s_weight7_bus_rreq_addr;
  -----------------------------------------------------------------------------
  s_weight0_bus_rdat_data                      <= s_bsv_rdat_data(BUS_DATA_WIDTH-1 downto 0);
  s_weight0_bus_rdat_last                      <= s_bsv_rdat_last(0);
  s_bsv_rdat_ready(0)                          <= s_weight0_bus_rdat_ready;
  s_weight0_bus_rdat_valid                     <= s_bsv_rdat_valid(0);
  -----------------------------------------------------------------------------
  s_weight1_bus_rdat_data                      <= s_bsv_rdat_data(2*BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH);
  s_bsv_rdat_ready(1)                          <= s_weight1_bus_rdat_ready;
  s_weight1_bus_rdat_valid                     <= s_bsv_rdat_valid(1);
  s_weight1_bus_rdat_last                      <= s_bsv_rdat_last(1);
  -----------------------------------------------------------------------------
  s_bsv_rdat_ready(2)                          <= s_weight2_bus_rdat_ready;
  s_weight2_bus_rdat_data                      <= s_bsv_rdat_data(3*BUS_DATA_WIDTH-1 downto 2*BUS_DATA_WIDTH);
  s_weight2_bus_rdat_last                      <= s_bsv_rdat_last(2);
  s_weight2_bus_rdat_valid                     <= s_bsv_rdat_valid(2);
  -----------------------------------------------------------------------------
  s_weight3_bus_rdat_valid                     <= s_bsv_rdat_valid(3);
  s_weight3_bus_rdat_last                      <= s_bsv_rdat_last(3);
  s_bsv_rdat_ready(3)                          <= s_weight3_bus_rdat_ready;
  s_weight3_bus_rdat_data                      <= s_bsv_rdat_data(4*BUS_DATA_WIDTH-1 downto 3*BUS_DATA_WIDTH);
  -----------------------------------------------------------------------------
  s_bsv_rdat_ready(4)                          <= s_weight4_bus_rdat_ready;
  s_weight4_bus_rdat_last                      <= s_bsv_rdat_last(4);
  s_weight4_bus_rdat_data                      <= s_bsv_rdat_data(5*BUS_DATA_WIDTH-1 downto 4*BUS_DATA_WIDTH);
  s_weight4_bus_rdat_valid                     <= s_bsv_rdat_valid(4);
  -----------------------------------------------------------------------------
  s_bsv_rdat_ready(5)                          <= s_weight5_bus_rdat_ready;
  s_weight5_bus_rdat_data                      <= s_bsv_rdat_data(6*BUS_DATA_WIDTH-1 downto 5*BUS_DATA_WIDTH);
  s_weight5_bus_rdat_last                      <= s_bsv_rdat_last(5);
  s_weight5_bus_rdat_valid                     <= s_bsv_rdat_valid(5);
  -----------------------------------------------------------------------------
  s_bsv_rdat_ready(6)                          <= s_weight6_bus_rdat_ready;
  s_weight6_bus_rdat_data                      <= s_bsv_rdat_data(7*BUS_DATA_WIDTH-1 downto 6*BUS_DATA_WIDTH);
  s_weight6_bus_rdat_valid                     <= s_bsv_rdat_valid(6);
  s_weight6_bus_rdat_last                      <= s_bsv_rdat_last(6);
  -----------------------------------------------------------------------------
  s_bsv_rdat_ready(7)                          <= s_weight7_bus_rdat_ready;
  s_weight7_bus_rdat_last                      <= s_bsv_rdat_last(7);
  s_weight7_bus_rdat_valid                     <= s_bsv_rdat_valid(7);
  s_weight7_bus_rdat_data                      <= s_bsv_rdat_data(8*BUS_DATA_WIDTH-1 downto 7*BUS_DATA_WIDTH);
  -----------------------------------------------------------------------------
  mst_wdat_valid                               <='0';
  mst_wreq_valid                               <='0';
  regs_out_en(0)                               <='0';
  regs_out_en(1)                               <='1';
  regs_out_en(2)                               <='1';
  regs_out_en(3)                               <='1';

end architecture;

